/*******************************************************************************************
*
*   raylib [textures] example - Load textures from raw data
*
*   NOTE: Images are loaded in CPU memory (RAM); textures are loaded in GPU memory (VRAM)
*
*   Example originally created with raylib 1.3, last time updated with raylib 3.5
*
*   Example licensed under an unmodified zlib/libpng license, which is an OSI-certified,
*   BSD-like license that allows static linking with closed source software
*
*   Copyright           (c) 2015-2023 Ramon Santamaria (@raysan5)
*   Translated&Modified (c) 2024      Fedorov Alexandr (@xydojnik)
*
********************************************************************************************/

module main


import raylib as rl


const asset_path  = @VMODROOT+'/thirdparty/raylib/examples/textures/resources/'


//------------------------------------------------------------------------------------
// Program main entry point
//------------------------------------------------------------------------------------
fn main() {
    // Initialization
    //--------------------------------------------------------------------------------------
    screen_width  := 800
    screen_height := 450

    rl.init_window(screen_width, screen_height, 'raylib [textures] example - texture from raw data')
    defer { rl.close_window() }                 // Close window and OpenGL context

    // NOTE: Textures MUST be loaded after Window initialization (OpenGL context is required)

    // Load RAW image data (512x512, 32bit RGBA, no file header)
    fudesumi_raw := rl.Image.load_raw(asset_path+'fudesumi.raw', 384, 512, rl.pixelformat_uncompressed_r8_g8_b8_a8, 0)
    fudesumi     := rl.load_texture_from_image(fudesumi_raw) // Upload CPU (RAM) image to GPU (VRAM)
    defer { fudesumi.unload() }                 // Texture unloading
    fudesumi_raw.unload()                       // Unload CPU (RAM) image data

    // Generate a checked texture by code
    mut width  := int(960)
    mut height := int(480)

    // Dynamic memory allocation to store pixels data (Color type)
    mut pixels := &rl.Color(rl.mem_alloc(u32(width*height)*sizeof(rl.Color)))

    for y in 0..height {
        for x in 0..width {
            unsafe {
                pixels[y*width+x] = if ((x/32+y/32)/1)%2 == 0 { rl.orange } else { rl.gold }
            }
        }
    }

    // Load pixels data into an image structure and create texture
    checked_im := rl.Image {
        data:     pixels,             // We can assign pixels directly to data
        width:    width,
        height:   height,
        format:   rl.pixelformat_uncompressed_r8_g8_b8_a8,
        mipmaps:  1
    }

    checked := rl.load_texture_from_image(checked_im)
    defer { rl.unload_texture(checked) } // Texture unloading
    rl.unload_image(checked_im)          // Unload CPU (RAM) image data (pixels)

    // Main game loop
    for !rl.window_should_close() {      // Detect window close button or ESC key
        // Update
        //----------------------------------------------------------------------------------
        // TODO: Update your variables here
        //----------------------------------------------------------------------------------

        // Draw
        //----------------------------------------------------------------------------------
        rl.begin_drawing()

            rl.clear_background(rl.raywhite)

            rl.draw_texture(checked, screen_width/2 - checked.width/2, screen_height/2 - checked.height/2, rl.Color.fade(rl.white, 0.5))
            rl.draw_texture(fudesumi, 430, -30, rl.white)

            rl.draw_text('CHECKED TEXTURE ',      84, 85 , 30, rl.brown)
            rl.draw_text('GENERATED by CODE',     72, 148, 30, rl.brown)
            rl.draw_text('and RAW IMAGE LOADING', 46, 210, 30, rl.brown)

            rl.draw_text('(c) Fudesumi sprite by Eiden Marsal', 310, screen_height - 20, 10, rl.brown)

        rl.end_drawing()
    }
}
