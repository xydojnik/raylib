module gui

#flag -DRAYGUI_IMPLEMENTATION

#include "@VMODROOT/../thirdparty/raylib/examples/shapes/raygui.h"
