module gui


pub const raygui_icon_size            = C.RAYGUI_ICON_SIZE             //  16  : Size of icons in pixels (squared)
pub const raygui_icon_max_icons       = C.RAYGUI_ICON_MAX_ICONS        //  256 : Maximum number of icons
pub const raygui_icon_max_name_length = C.RAYGUI_ICON_MAX_NAME_LENGTH  //  32  : Maximum length of icon name id

pub const raygui_icon_data_elements   = C.RAYGUI_ICON_DATA_ELEMENTS

pub const gui_icons                   = C.guiIcons

pub const scrollbar_left_side         = C.SCROLLBAR_LEFT_SIDE   // 0
pub const scrollbar_right_side        = C.SCROLLBAR_RIGHT_SIDE  // 1
