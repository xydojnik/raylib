module gui

#flag -DRAYGUI_IMPLEMENTATION

#include "@VMODROOT/raygui.h"
